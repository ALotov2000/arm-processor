module ControlUnit(
    input[3:0] opcode, 
    input[1:0] mode, 
    input S_in, 

    output[8:0] out
);

endmodule